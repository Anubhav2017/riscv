module data_mem(
    input [4:0] rdaddr1, rdaddr2, wraddr1
);


endmodule
module riscv_top();



endmodule